Library ieee;
use ieee.std_logic_1164.all;
use work.Comp_package.all;
entity MIPS is
	port(	 
		 rst : in std_logic
		);	  
end MIPS;


architecture arch of MIPS is
signal pcOut :  std_logic_vector(31 downto 0);
signal instruct_memory : std_logic_vector(31 downto 0);
signal outControlUnit : std_logic_vector(12 downto 0);
signal pcAdderOut : std_logic_vector(31 downto 0);
signal outmux1: std_logic_vector(4 downto 0); 
signal outmux32bit2: std_logic_vector(31 downto 0);
signal readdata1: std_logic_vector(31 downto 0);
signal readdata2: std_logic_vector(31 downto 0);	 
signal ot_si_ex : std_logic_vector(31 downto 0); 
signal outmux32bit1: std_logic_vector(31 downto 0); 
signal out_alu_control: std_logic_vector(5 downto 0);
signal zero : STD_LOGIC;							 
signal alu_result : std_logic_vector(31 downto 0);	
signal datamemory_out : std_logic_vector(31 downto 0); 
signal shiftleftout2: std_logic_vector(31 downto 0); 
signal addout: std_logic_vector(31 downto 0);
signal outmux32bit3: std_logic_vector(31 downto 0);	
signal outandgate: std_logic;  
 signal clk1,clk2,clk3,clk4: std_logic:='1';	--1-pc   2- regread 3- regwrite 4 -dm 
begin
	
	process is
    begin 
		while(true) loop
        clk1 <= not clk1;  
		wait for 200 ps;
		end loop;
    end process;

    process is
    begin 
        wait for 50 ps;
        while(true) loop
            clk2 <= not clk2;
            wait for 200 ps;
        end loop; 
    end process;

    process is
    begin	  
        wait for 100 ps;
        while(true) loop
            clk4 <= not clk4;
            wait for 200 ps;
        end loop;
    end process;

    process is
	begin  
            wait for 150 ps;
            while(true) loop
                clk3 <= not clk3;
                wait for 200 ps;
            end loop;
    end process;


	pc : entity work.ProgramCounter port map  (clk1,rst,outmux32bit3 ,pcOut);
	insmemory : entity work.InstructionMemory port map(clk1,pcOut, instruct_memory);
	CU :  entity work.ControlUnit port map(instruct_memory(31 downto 26),
	outControlUnit(0),  
	outControlUnit(1),
	outControlUnit(2),
	outControlUnit(3),
	outControlUnit(4),
	outControlUnit(5),
	outControlUnit(6),
	outControlUnit(12 downto 7));
	
	muxinstructionmemroytoregister: entity work.mux5bit port map(instruct_memory(20 downto 16),
	instruct_memory(15 downto 11), outControlUnit(0),outmux1); 
	
	pcAdder : entity work.ProgramCounterAdder port map(pcOut, pcAdderOut); 
	
	reg_file : entity work.RegisterFile port map(clk2,clk3,outControlUnit(3),outmux1, outmux32bit2,
	instruct_memory(25 downto 21),instruct_memory(20 downto 16), readdata1, readdata2);
	
	sign : entity work.SignExtender port map  (instruct_memory(15 downto 0) ,ot_si_ex);
	
	mux32bit: entity work.MUX port map(readdata2,ot_si_ex,outControlUnit(1),outmux32bit1);
	
	alu  : entity work.ALU port map (out_alu_control,readdata1,outmux32bit1,alu_result,zero); 
	alu_control : entity work.ALU_Control port map (instruct_memory(5 downto 0),
	outControlUnit(12 downto 7) ,out_alu_control) ;		 
	
	datamemorylabel : entity work.DataMemory port map ( clk4,alu_result,
	readdata2,outControlUnit(4),outControlUnit(5), datamemory_out);	
	
	mux32bit2 : entity work.MUX port map(alu_result,datamemory_out,outControlUnit(2),outmux32bit2);	 
	shiftL1 : entity work.Shift2Left port map(ot_si_ex, shiftleftout2);	
	
	adder: entity work.adder port map(pcAdderOut,shiftleftout2, addout);	  
	
	mux32bit3 : entity work.MUX port map(pcAdderOut,addout, outandgate,outmux32bit3);  
	andgate: entity work.andgate port map(zero,outControlUnit(6), outandgate); 
end arch;